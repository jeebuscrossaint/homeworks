library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Mux16to1_AmarnathPatelVHDL is
    Port(
        sel : in STD_LOGIC_VECTOR(3 downto 0);  -- 4 selection bits
        in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11,in12,in13,in14,in15  : in STD_LOGIC;  -- Input 0
        output : out STD_LOGIC -- Output
    );
end Mux16to1_AmarnathPatelVHDL;

architecture structural of Mux16to1_AmarnathPatelVHDL is
    -- Component declarations
    component Mux4to1_AmarnathPatelVHDL is
        Port(
            sel : in STD_LOGIC_VECTOR(1 downto 0);
            in0, in1, in2, in3 : in STD_LOGIC;
            output : out STD_LOGIC
        );
    end component;
    
    component Mux2to1_AmarnathPatelVHDL is
        Port(
            s,x,y : in STD_LOGIC;
 
            mux : out STD_LOGIC
        );
    end component;
    
    -- Internal signals for intermediate MUX outputs
    signal mux4to1_out1 : STD_LOGIC;  -- Output from first 4:1 MUX
    signal mux4to1_out2 : STD_LOGIC;  -- Output from second 4:1 MUX
    signal mux4to1_out3 : STD_LOGIC;  -- Output from third 4:1 MUX
    signal mux4to1_out4 : STD_LOGIC;  -- Output from fourth 4:1 MUX
    signal mux2to1_out1 : STD_LOGIC;  -- Output from first 2:1 MUX
    signal mux2to1_out2 : STD_LOGIC;  -- Output from second 2:1 MUX
    
begin
    -- First level: Four 4-to-1 MUXes
    MUX4_1: Mux4to1_AmarnathPatelVHDL
        port map(
            sel => sel(1 downto 0),
            in0 => in0,
            in1 => in1,
            in2 => in2,
            in3 => in3,
            output => mux4to1_out1
        );
        
    MUX4_2: Mux4to1_AmarnathPatelVHDL
        port map(
            sel => sel(1 downto 0),
            in0 => in4,
            in1 => in5,
            in2 => in6,
            in3 => in7,
            output => mux4to1_out2
        );
        
    MUX4_3: Mux4to1_AmarnathPatelVHDL
        port map(
            sel => sel(1 downto 0),
            in0 => in8,
            in1 => in9,
            in2 => in10,
            in3 => in11,
            output => mux4to1_out3
        );
        
    MUX4_4: Mux4to1_AmarnathPatelVHDL
        port map(
            sel => sel(1 downto 0),
            in0 => in12,
            in1 => in13,
            in2 => in14,
            in3 => in15,
            output => mux4to1_out4
        );
        
    -- Second level: Two 2-to-1 MUXes
    MUX2_1: Mux2to1_AmarnathPatelVHDL
        port map(
            s => sel(2),
            x => mux4to1_out1,
            y => mux4to1_out2,
            mux => mux2to1_out1
        );
        
    MUX2_2: Mux2to1_AmarnathPatelVHDL
        port map(
            s => sel(2),
            x => mux4to1_out3,
            y => mux4to1_out4,
            mux => mux2to1_out2
        );
        
    -- Final level: One 2-to-1 MUX
    MUX2_FINAL: Mux2to1_AmarnathPatelVHDL
        port map(
            s => sel(3),
            x => mux2to1_out1,
            y => mux2to1_out2,
            mux => output
        );
        
end structural;