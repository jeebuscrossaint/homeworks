LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;

ENTITY NAND4_AmarnathPatelVHDL is
	PORT(X0,X1,X2,X3:IN STD_LOGIC;
					:OUT STD_LOGIC);
END NAND4_AmarnathPatelVHDL;

ARCHITECTURE Structure OF NAND4_AmarnathPatelVHDL is
BEGIN

f <=(((X0 NAND X1) NAND (X0 NAND X1))NAND((X2 NAND X3)NAND(X2 NAND X3)));

END Structure