LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;

ENTITY NAND3_AmarnathPatelVHDL is
	PORT(X0,X1,X2:IN STD_LOGIC;
		 f		 :OUT STD_LOGIC);
END NAND3_AmarnathPatelVHDL;

ARCHITECTURE Structure OF NAND3_AmarnathPatelVHDL IS
BEGIN

f <= (((X0 NAND X1)NAND(X0 NAND X1))NAND X2);

END Structure